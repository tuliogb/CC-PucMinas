/*
	Nome: Tulio Gomes Braga 
	Matricula: 802512	
*/

`include "clock.v"

module pulse1 ( signal, clock );
    input clock;
    output signal;
    reg signal;
    
    always @ ( posedge clock ) begin
        signal = 1'b1;
        #2 signal = 1'b0;
        #2 signal = 1'b1;
        #2 signal = 1'b0;
        #2 signal = 1'b1;
        #2 signal = 1'b0;
    end
endmodule

module Guia_0905;
    wire clock;
    clock clk ( clock );
    wire p1;

    pulse1 pls1( p1, clock );

    initial begin
        $dumpfile ( "Guia_0905.vcd" );
        $dumpvars ( 1, clock, p1);	
        #240 $finish;
    end
endmodule 


/*
	Se o clock estiver em borda de subida(1), de 2 em 2 segundo sao gerados pulsos.
*/
